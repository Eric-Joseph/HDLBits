module top_module(
    input clk,
    input a,
    input b,
    output wire out_assign,
    output reg out_always_comb,
    output reg out_always_ff   );

endmodule

// UNDER DEVELOPMENT. WILL FINISH AT A LATER DATE
